module psi

pub interface PsiDocCommentOwner {
	doc_comment() string
}
