module psi

pub struct PlainType {
	PsiElementImpl
}

fn (_ &PlainType) stub() {}
