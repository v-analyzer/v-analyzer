// MIT License
//
// Copyright (c) 2023-2024 V Open Source Community Association (VOSCA) vosca.dev
//
// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:
//
// The above copyright notice and this permission notice shall be included in all
// copies or substantial portions of the Software.
//
// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
// SOFTWARE.
module stubs

// err is a special variable that is set with an error
// and is used to handle errors in V.
//
// It can be used inside two places:
//
// 1. inside `or` block:
// ```
// fn foo() !int {
//   return error("not implemented");
// }
//
// foo() or {
//   panic(err);
//   //    ^^^ err is set with error("not implemented")
// }
// ```
//
// 2. inside else block for if guard:
// ```
// fn foo() !int {
//   return error("not implemented");
// }
//
// if val := foo() {
//   // val is set with int
// } else {
//   panic(err);
//   //    ^^^ err is set with error("not implemented")
// }
// ```
//
// See [Documentation](https://docs.vosca.dev/concepts/error-handling/overview.html)
// for more details.
pub const err = IError{}
