module types

struct BaseType {
}
