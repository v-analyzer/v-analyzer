module psi

pub struct Argument {
	PsiElementImpl
}
