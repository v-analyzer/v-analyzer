module psi

pub interface SignatureOwner {
	signature() ?&Signature
}
