// MIT License
//
// Copyright (c) 2023-2024 V Open Source Community Association (VOSCA) vosca.dev
//
// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:
//
// The above copyright notice and this permission notice shall be included in all
// copies or substantial portions of the Software.
//
// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
// SOFTWARE.
module main

import testing

fn bench() testing.BenchmarkRunner {
	mut b := testing.BenchmarkRunner{
		last_fixture: unsafe { nil }
	}

	b.bench('inlay hints', fn (mut b testing.Benchmark, mut fixture testing.Fixture) ! {
		fixture.configure_by_file('benchmarks/checker.v')!

		b.start()

		hints := fixture.compute_inlay_hints()
		println('Count: ${hints.len}')

		b.stop()
		b.print_results()
	})

	b.bench('semantic tokens', fn (mut b testing.Benchmark, mut fixture testing.Fixture) ! {
		fixture.configure_by_file('benchmarks/checker.v')!

		b.start()

		tokens := fixture.compute_semantic_tokens()
		println('Count: ${tokens.data.len / 5}')

		b.stop()
		b.print_results()
	})

	return b
}
