module indexer

pub struct PerFileCache {
pub mut:
	data map[string]Cache
}
