module types

struct FooBar {
}

fn some_foo() string {}

fn foo_int() int {}

fn get_foo_bar() FooBar {}

fn main() {
	expr_type(some_foo(), 'string')
	expr_type(foo_int(), 'int')
	expr_type(get_foo_bar(), 'types.FooBar')
}
