module indexer

// Index инкапсулирует логику хранения индекса.
pub struct Index {
	version string = '0.0.1'
}
