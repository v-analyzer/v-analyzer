module psi

pub struct ParameterList {
	PsiElementImpl
}

fn (n &ParameterList) stub() {}
