module psi

pub struct Signature {
	PsiElementImpl
}
