module types

fn main() {
	expr_type(100, 'int')
	expr_type(3.14, 'f64')
	expr_type(`r`, 'rune')
	expr_type(true, 'bool')
	expr_type(false, 'bool')
	expr_type(nil, 'voidptr')
	expr_type(none, 'none')
	expr_type('hello', 'string')
	expr_type(r'raw hello', 'string')
	expr_type(c'c hello', '&u8')
}
