module psi

pub struct Comment {
	PsiElementImpl
}
