// MIT License
//
// Copyright (c) 2023-2024 V Open Source Community Association (VOSCA) vosca.dev
//
// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:
//
// The above copyright notice and this permission notice shall be included in all
// copies or substantial portions of the Software.
//
// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
// SOFTWARE.
module server

import lsp
import loglib

pub fn (mut ls LanguageServer) did_change_watched_files(params lsp.DidChangeWatchedFilesParams) {
	changes := params.changes
	mut is_rename := false

	// NOTE:
	// 1. Renaming a file returns two events: one "created" event for the
	//    same file with new name and one "deleted" event for the file with
	//    old name.
	// 2. Deleting a folder does not trigger a "deleted" event. Restoring
	//    the files of the folder however triggers the "created" event.
	// 3. Renaming a folder triggers the "created" event for each file
	//    but with no "deleted" event prior to it.
	for i, change in changes {
		change_uri := change.uri.normalize()
		match change.typ {
			.created {
				if next_change := changes[i + 1] {
					is_rename = next_change.typ == .deleted
				}

				if is_rename {
					prev_change := changes[i + 1] or { continue }
					prev_uri := prev_change.uri.normalize()
					if file_index := ls.indexing_mng.indexer.rename_file(prev_uri.path(),
						change_uri.path())
					{
						if isnil(file_index.sink) {
							continue
						}

						ls.indexing_mng.update_stub_indexes_from_sinks([*file_index.sink])

						loglib.with_fields({
							'old': prev_uri.path()
							'new': change_uri.path()
						}).info('Renamed file')
					}
				} else {
					if file_index := ls.indexing_mng.indexer.add_file(change_uri.path()) {
						if isnil(file_index.sink) {
							continue
						}

						ls.indexing_mng.update_stub_indexes_from_sinks([*file_index.sink])

						loglib.with_fields({
							'file': change_uri.path()
						}).info('Added file')
					}
				}
			}
			.deleted {
				if is_rename {
					continue
				}
				if file_index := ls.indexing_mng.indexer.remove_file(change_uri.path()) {
					if isnil(file_index.sink) {
						continue
					}

					ls.indexing_mng.update_stub_indexes_from_sinks([*file_index.sink])

					loglib.with_fields({
						'file': change_uri.path()
					}).info('Removed file')
				}
			}
			.changed {}
		}

		ls.client.log_message(change.str(), .info)
	}
}
