module psi

pub struct ImportName {
	PsiElementImpl
}

fn (n &ImportName) stub() {}
