module psi

pub struct ImportDeclaration {
	PsiElementImpl
}

fn (n &ImportDeclaration) stub() {}
