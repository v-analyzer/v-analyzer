module psi

pub interface PsiComment {
	PsiElement
	get_content() string
}
