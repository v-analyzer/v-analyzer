module psi

pub interface AttributesOwner {
	attributes() []Attribute
}
