module psi

pub interface AttributesOwner {
	attributes() []PsiElement
}
