module psi

pub struct Position {
pub:
	line      int
	character int
}
