// MIT License
//
// Copyright (c) 2023-2024 V Open Source Community Association (VOSCA) vosca.dev
//
// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:
//
// The above copyright notice and this permission notice shall be included in all
// copies or substantial portions of the Software.
//
// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
// SOFTWARE.
module lsp

// method: ‘textDocument/formatting’
// response: []TextEdit | none
pub struct DocumentFormattingParams {
pub:
	text_document TextDocumentIdentifier @[json: textDocument]
	options       FormattingOptions
}

pub struct FormattingOptions {
	tab_size      int  @[json: tabSize]
	insert_spaces bool @[json: insertSpaces]
	// [key] bool | number | string
}

// method: ‘textDocument/rangeFormatting’
// response: []TextEdit | none
pub struct DocumentRangeFormattingParams {
	text_document TextDocumentIdentifier @[json: textDocument]
	range         Range
	options       FormattingOptions
}

pub struct DocumentOnTypeFormattingOptions {
	first_trigger_character string   @[json: firstTriggerCharacter]
	more_trigger_character  []string @[json: moreTriggerCharacter]
}

// method: ‘textDocument/onTypeFormatting’
// response: []TextEdit | none
pub struct DocumentOnTypeFormattingParams {
	text_document TextDocumentIdentifier @[json: textDocument]
	position      Position
	ch            string
	options       FormattingOptions
}

pub struct DocumentOnTypeFormattingRegistrationOptions {
	document_selector       []DocumentFilter @[json: documentSelector]
	first_trigger_character string           @[json: firstTriggerCharacter]
	more_trigger_character  []string         @[json: moreTriggerCharacter]
}
