module main

import net.http

type Foo = string

struct Goo {}

fn foo() {
	name, some, mut other := "", 1, 2

	println(name)
	println(some)
	println(other)

	if 1 {
		name := 11
		println(name)
		println(some)
	}
}

foo()
Foo
	Goo{}

foo.goo.zoo
http.foo()


