module psi

[heap]
pub struct StubIndexSink {
pub mut:
	stub_id     StubId
	stub_list   &StubList // Список стаблв в текущем файле для которого строится индекс
	module_name string
	data        map[int]map[string][]StubId
}

fn (mut s StubIndexSink) occurrence(key StubIndexKey, value string) {
	resulting_value := if s.module_name != '' {
		s.module_name + '.' + value
	} else {
		value
	}

	mut values := s.data[int(key)].move()
	values[resulting_value] << s.stub_id
	s.data[int(key)] = values.move()
}
