module psi

pub interface GenericParametersOwner {
	generic_parameters() ?&GenericParameters
}
