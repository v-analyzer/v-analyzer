module types

fn main() {
	a := 100
	expr_type(a, 'int')
}
