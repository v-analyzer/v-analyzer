module psi

pub struct ImportAlias {
	PsiElementImpl
}

fn (n &ImportAlias) stub() {}
