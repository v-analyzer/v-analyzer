// MIT License
//
// Copyright (c) 2023-2024 V Open Source Community Association (VOSCA) vosca.dev
//
// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:
//
// The above copyright notice and this permission notice shall be included in all
// copies or substantial portions of the Software.
//
// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
// SOFTWARE.
module attributes

// JsonAsNumber marks an enum.
// The fields of such enum will be encoded in JSON as numbers, not as strings
// with the field name.
//
// Example:
//
// ```
// [json_as_number]
// enum Color {
//   red = 1
//   green = 2
// }
//
// struct MyStruct {
//   color Color = .green
// }
//
// // JSON representation of MyStruct:
// // {
// //   "color": 2
// // }
//
// // JSON representation of MyStruct without the attribute:
// // {
// //   "color": "green"
// // }
// ```
@[attribute]
pub struct JsonAsNumber {
	name            string = 'json_as_number'
	with_arg        bool
	arg_is_optional bool
	target          []Target = [Target.enum_]
}
