module types

fn main() {
	ch := chan int{}
	expr_type(ch, 'chan int')
	expr_type(<-ch, 'int')
}
