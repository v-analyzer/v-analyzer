// MIT License
//
// Copyright (c) 2023-2024 V Open Source Community Association (VOSCA) vosca.dev
//
// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:
//
// The above copyright notice and this permission notice shall be included in all
// copies or substantial portions of the Software.
//
// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
// SOFTWARE.
module lsp

pub struct CodeLensOptions {
pub mut:
	resolve_provider   bool @[json: 'resolveProvider'; omitempty]
	work_done_progress bool @[json: 'workDoneProgress'; omitempty]
}

// method: ‘textDocument/codeLens’
// response: []CodeLens | none
pub struct CodeLensParams {
	WorkDoneProgressParams
pub:
	text_document TextDocumentIdentifier @[json: textDocument]
}

pub struct CodeLens {
pub:
	// The range in which this code lens is valid. Should only span a single
	// line.
	range Range
	// The command this code lens represents.
	command Command
	// A data entry field that is preserved on a code lens item between
	// a code lens and a code lens resolve request.
	data string @[raw]
}

pub struct CodeLensRegistrationOptions {
	document_selector []DocumentFilter @[json: documentSelector]
	resolve_provider  bool             @[json: resolveProvider]
}

// method: ‘codeLens/resolve’
// response: CodeLens
// request: CodeLens
