module types

fn main() {
	a := 100
	b := &a
	c := &b
	d := *c
	e := *d

	expr_type(a, 'int')
	expr_type(b, '&int')
	expr_type(c, '&&int')
	expr_type(d, '&int')
	expr_type(e, 'int')
}
