module documentation

// has checks if the enum value has the passed flag.
//
// **bold**
// *italic*
// `code`
// [link](https://github.com)
// ---
//
// # Heading 1
// ## Heading 2
// ### Heading 3
//
// line break.
// line break!
// line break?
//
// Example:
// ```
// [flag]
// enum Permissions {
//   read  // = 0b0001
//   write // = 0b0010
//   other // = 0b0100
// }
//
// fn main() {
//   p := Permissions.read
//   assert p.has(.read) // test if p has read flag
//   assert p.has(.read | .other) // test if *at least one* of the flags is set
// }
// ```
//
// Example: println('inline example')
fn foo() { // caret
}
