module psi

pub struct FieldName {
	PsiElementImpl
}
