module psi

pub struct ParameterList {
	PsiElementImpl
}

fn (_ &ParameterList) stub() {}
