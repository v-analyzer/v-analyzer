module psi

pub struct ImportList {
	PsiElementImpl
}

fn (n &ImportList) stub() {}
