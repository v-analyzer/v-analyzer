module psi

pub struct TextRange {
pub:
	line       int
	column     int
	end_line   int
	end_column int
}
