// MIT License
//
// Copyright (c) 2023-2024 V Open Source Community Association (VOSCA) vosca.dev
//
// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:
//
// The above copyright notice and this permission notice shall be included in all
// copies or substantial portions of the Software.
//
// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
// SOFTWARE.
module attributes

// Noreturn attribute marks a function as not return to its caller.
//
// Such functions can be used at the end of or blocks, just like
// [`exit`](#exit) or [`panic`](#panic).
//
// Such functions can not have return types, and should end either in `for {}`, or
// by calling other `[noreturn]` functions.
//
// Example:
//
// ```
// [noreturn]
// fn redirect() {
//    // do something
//    exit(1)
// }
//
// fn main() {
//     if condition {
//         redirect();
//         // unreachable
//     }
// }
// ```
@[attribute]
pub struct Noreturn {
	name            string = 'noreturn'
	with_arg        bool
	arg_is_optional bool
	target          []Target = [Target.function]
}
