module types

expr_type(unsafe { 100 }, 'int')
expr_type(unsafe {
	a := 100
	a
}, 'int')
