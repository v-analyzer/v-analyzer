// MIT License
//
// Copyright (c) 2023-2024 V Open Source Community Association (VOSCA) vosca.dev
//
// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:
//
// The above copyright notice and this permission notice shall be included in all
// copies or substantial portions of the Software.
//
// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
// SOFTWARE.
module types

fn main() {
	a := if true {
		100
	} else {
		200
	}
	expr_type(a, 'int')

	b := if true {
		'100'
	} else {
		'200'
	}
	expr_type(b, 'string')

	c := if true {
		unsafe { 100 }
	} else {
		200
	}
	expr_type(c, 'int')

	d := if true {
		inner := unsafe { 100 }
		inner
	} else {
		200
	}
	expr_type(d, 'int')

	e := if true {
		inner := map[int]string{}
		inner[100]
	} else {
		200
	}
	expr_type(e, 'string')

	f := if true {
		unknown
	} else {
		200
	}
	expr_type(f, 'int')

	g := $if macos {
		1
	} $else {
		2
	}
	expr_type(g, 'int')
}

fn get_opt() ?int {
	return 100
}

fn get_res() !int {
	return 100
}

fn unwrapping() {
	if a := get_opt() {
		expr_type(a, 'int')
	}

	if a := get_res() {
		expr_type(a, 'int')
	}
}
