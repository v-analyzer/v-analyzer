module types

struct ReceiverFoo {}

fn (r &ReceiverFoo) method() {
	expr_type(r, '&types.ReceiverFoo')
	expr_type(*r, 'types.ReceiverFoo')
}
