module psi

@[heap]
pub struct PlainType {
	PsiElementImpl
}

fn (_ &PlainType) stub() {}
