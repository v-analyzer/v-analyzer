module psi

pub struct ImportPath {
	PsiElementImpl
}

fn (n &ImportPath) stub() {}
