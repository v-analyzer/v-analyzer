module psi

pub struct MutExpression {
	PsiElementImpl
}
