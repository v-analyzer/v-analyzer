module psi

// StubIndexKey описывает различные типы индексов, которые строятся
// по `index.StubTree`.
// Эти индексы позволяют быстро находить нужные определения по имени
// во всех проиндексированных файлах, включая стандартную библиотеку и
// сторонние библиотеки вне проекта.
pub enum StubIndexKey as u8 {
	functions
	methods
	structs
	constants
	type_aliases
	enums
	attributes
}

// IndexSink описывает интерфейс создателя индексов.
// Метод `occurrence()` вызывается для каждого стаба в файле. Смотри
// `StubbedElementType.index_stub()` для примера вызова этого метода.
//
// Параметр `key` это тип индекса, для которого нужно создать запись.
// Параметр `value` это строка, которая будет использована в качестве
// значения в индексе. Например, для индекса `functions` это будет имя функции.
pub interface IndexSink {
mut:
	occurrence(key StubIndexKey, value string)
}

// StubBasedPsiElement описывает маркерный интерфейс для элементов PSI,
// из которых будет построено `index.StubTree`, по которому будут построены
// стабовые индексы.
//
// PSI элементы которые реализуют этот интерфейс могут быть созданы
// как из AST, так и из стабов (`psi.StubBase`).
// Это позволяет единообразно обрабатывать их при резолвинге имен и
// другой обработке, так как нет разницы, обрабатываем мы реальное AST
// дерево или дерево стабов из память.
pub interface StubBasedPsiElement {
	stub() // marker method
}
