module psi

pub struct ParameterDeclaration {
	PsiElementImpl
}
