// MIT License
//
// Copyright (c) 2023-2024 V Open Source Community Association (VOSCA) vosca.dev
//
// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:
//
// The above copyright notice and this permission notice shall be included in all
// copies or substantial portions of the Software.
//
// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
// SOFTWARE.
module types

fn arrays() {
	for index in 0 .. 10 {
		expr_type(index, 'int')
	}

	int_array := [1, 2, 3]

	for index in int_array {
		expr_type(index, 'int')
	}

	for index, value in int_array {
		expr_type(index, 'int')
		expr_type(value, 'int')
	}

	string_array := ['1', '2', '3']

	for index in string_array {
		expr_type(index, 'string')
	}

	for index, value in string_array {
		expr_type(index, 'int')
		expr_type(value, 'string')
	}

	bool_array := [true, false]

	for index in bool_array {
		expr_type(index, 'bool')
	}

	for index, value in bool_array {
		expr_type(index, 'int')
		expr_type(value, 'bool')
	}
}

fn maps() {
	mp := map[string]int{}

	for key, value in mp {
		expr_type(key, 'string')
		expr_type(value, 'int')
	}
}

fn strings() {
	mp := ''

	for value in mp {
		expr_type(value, 'u8')
	}

	for key, value in mp {
		expr_type(key, 'int')
		expr_type(value, 'u8')
	}
}
